`define WIDTH 7
