`define WIDTH 7
`define NUM_CANDIDATES 3
`define MAX_WAIT_CYCLE 101
