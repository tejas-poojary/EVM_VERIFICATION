`define WIDTH 7
`define NUM_CANDIDATES 3
