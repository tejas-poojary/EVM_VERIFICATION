package evm_pkg;
`include "evm_sequence_item.sv"
`include "evm_sequence.sv"
`include "evm_sequencer.sv"
`include "evm_driver.sv"
`include "evm_active_monitor.sv"
`include "evm_passive_monitor.sv"
`include "evm_agent.sv"
`include "evm_scoreboard.sv"
`include "evm_subscriber.sv"
`include "evm_environment.sv"
`include "evm_test.sv"
endpackage
